MACRO Bimod_Tag_ROM
  PIN A[0]
    ANTENNAGATEAREA 0.0224 ;
    ANTENNADIFFAREA 0.096 ;
    END A[0]
  PIN A[1]
    ANTENNAGATEAREA 0.0224 ;
    ANTENNADIFFAREA 0.096 ;
    END A[1]
  PIN A[2]
    ANTENNAGATEAREA 0.0224 ;
    ANTENNADIFFAREA 0.096 ;
    END A[2]
  PIN A[3]
    ANTENNAGATEAREA 0.0224 ;
    ANTENNADIFFAREA 0.096 ;
    END A[3]
  PIN A[4]
    ANTENNAGATEAREA 0.0224 ;
    ANTENNADIFFAREA 0.096 ;
    END A[4]
  PIN A[5]
    ANTENNAGATEAREA 0.0224 ;
    ANTENNADIFFAREA 0.096 ;
    END A[5]
  PIN A[6]
    ANTENNAGATEAREA 0.0224 ;
    ANTENNADIFFAREA 0.096 ;
    END A[6]
  PIN CEN
    ANTENNAGATEAREA 0.0224 ;
    ANTENNADIFFAREA 0.096 ;
    END CEN
  PIN CLK
    ANTENNAGATEAREA 0.0224 ;
    ANTENNADIFFAREA 0.096 ;
    END CLK
  END Bimod_Tag_ROM ;
  END LIBRARY
