library verilog;
use verilog.vl_types.all;
entity test_top is
end test_top;
